library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;
use ieee.numeric_std.all;

package arr_package is

	type input_arr is array(0 to 10) of std_logic_vector(47 downto 0); 
	type output_arr is array(0 to 10) of std_logic_vector(7 downto 0); 
  
end package arr_package;
 
-- Package Body Section
package body arr_package is
 

 
end package body arr_package;